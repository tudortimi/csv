module automatic dict_writer_example;
    import csv::*;
endmodule
